module dut();
  initial 
    $hello();
endmodule // test